#
# Automatically generated make config: don't edit
# Busybox version: 1.36.0
# Fri Jan 27 09:01:31 2023
#
CONFIG_HAVE_DOT_CONFIG=y

#
# Settings
#
# CONFIG_DESKTOP is not set
# CONFIG_EXTRA_COMPAT is not set
# CONFIG_FEDORA_COMPAT is not set
# CONFIG_INCLUDE_SUSv2 is not set
CONFIG_LONG_OPTS=y
CONFIG_SHOW_USAGE=y
CONFIG_FEATURE_VERBOSE_USAGE=y
CONFIG_FEATURE_COMPRESS_USAGE=y
# CONFIG_LFS is not set
# CONFIG_PAM is not set
# CONFIG_FEATURE_DEVPTS is not set
# CONFIG_FEATURE_UTMP is not set
# CONFIG_FEATURE_WTMP is not set
# CONFIG_FEATURE_PIDFILE is not set
CONFIG_PID_FILE_PATH=""
CONFIG_BUSYBOX=y
CONFIG_FEATURE_SHOW_SCRIPT=y
CONFIG_FEATURE_INSTALLER=y
CONFIG_INSTALL_NO_USR=y
# CONFIG_FEATURE_SUID is not set
# CONFIG_FEATURE_SUID_CONFIG is not set
# CONFIG_FEATURE_SUID_CONFIG_QUIET is not set
# CONFIG_FEATURE_PREFER_APPLETS is not set
CONFIG_BUSYBOX_EXEC_PATH="/proc/self/exe"
# CONFIG_SELINUX is not set
# CONFIG_FEATURE_CLEAN_UP is not set
CONFIG_FEATURE_SYSLOG_INFO=y
CONFIG_FEATURE_SYSLOG=y

#
# Build Options
#
CONFIG_STATIC=y
# CONFIG_PIE is not set
# CONFIG_NOMMU is not set
# CONFIG_BUILD_LIBBUSYBOX is not set
# CONFIG_FEATURE_LIBBUSYBOX_STATIC is not set
# CONFIG_FEATURE_INDIVIDUAL is not set
# CONFIG_FEATURE_SHARED_BUSYBOX is not set
CONFIG_CROSS_COMPILER_PREFIX="x86_64-linux-android-"
CONFIG_SYSROOT=""
CONFIG_EXTRA_CFLAGS=""
CONFIG_EXTRA_LDFLAGS=""
CONFIG_EXTRA_LDLIBS=""
# CONFIG_USE_PORTABLE_CODE is not set
CONFIG_STACK_OPTIMIZATION_386=y
CONFIG_STATIC_LIBGCC=y

#
# Installation Options ("make install" behavior)
#
CONFIG_INSTALL_APPLET_SYMLINKS=y
# CONFIG_INSTALL_APPLET_HARDLINKS is not set
# CONFIG_INSTALL_APPLET_SCRIPT_WRAPPERS is not set
# CONFIG_INSTALL_APPLET_DONT is not set
# CONFIG_INSTALL_SH_APPLET_SYMLINK is not set
# CONFIG_INSTALL_SH_APPLET_HARDLINK is not set
# CONFIG_INSTALL_SH_APPLET_SCRIPT_WRAPPER is not set
CONFIG_PREFIX="./_install"

#
# Debugging Options
#
# CONFIG_DEBUG is not set
# CONFIG_DEBUG_PESSIMIZE is not set
# CONFIG_DEBUG_SANITIZE is not set
# CONFIG_UNIT_TEST is not set
# CONFIG_WERROR is not set
# CONFIG_WARN_SIMPLE_MSG is not set
CONFIG_NO_DEBUG_LIB=y
# CONFIG_DMALLOC is not set
# CONFIG_EFENCE is not set

#
# Library Tuning
#
# CONFIG_FEATURE_USE_BSS_TAIL is not set
CONFIG_FLOAT_DURATION=y
# CONFIG_FEATURE_RTMINMAX is not set
# CONFIG_FEATURE_RTMINMAX_USE_LIBC_DEFINITIONS is not set
CONFIG_FEATURE_BUFFERS_USE_MALLOC=y
# CONFIG_FEATURE_BUFFERS_GO_ON_STACK is not set
# CONFIG_FEATURE_BUFFERS_GO_IN_BSS is not set
CONFIG_PASSWORD_MINLEN=6
CONFIG_MD5_SMALL=1
CONFIG_SHA1_SMALL=3
CONFIG_SHA1_HWACCEL=y
CONFIG_SHA256_HWACCEL=y
CONFIG_SHA3_SMALL=1
# CONFIG_FEATURE_NON_POSIX_CP is not set
CONFIG_FEATURE_VERBOSE_CP_MESSAGE=y
CONFIG_FEATURE_USE_SENDFILE=y
CONFIG_FEATURE_COPYBUF_KB=4
# CONFIG_MONOTONIC_SYSCALL is not set
# CONFIG_IOCTL_HEX2STR_ERROR is not set
CONFIG_FEATURE_EDITING=y
CONFIG_FEATURE_EDITING_MAX_LEN=1024
CONFIG_FEATURE_EDITING_VI=y
CONFIG_FEATURE_EDITING_HISTORY=255
CONFIG_FEATURE_EDITING_SAVEHISTORY=y
# CONFIG_FEATURE_EDITING_SAVE_ON_EXIT is not set
CONFIG_FEATURE_REVERSE_SEARCH=y
CONFIG_FEATURE_TAB_COMPLETION=y
# CONFIG_FEATURE_USERNAME_COMPLETION is not set
CONFIG_FEATURE_EDITING_FANCY_PROMPT=y
CONFIG_FEATURE_EDITING_WINCH=y
# CONFIG_FEATURE_EDITING_ASK_TERMINAL is not set
# CONFIG_LOCALE_SUPPORT is not set
# CONFIG_UNICODE_SUPPORT is not set
# CONFIG_UNICODE_USING_LOCALE is not set
# CONFIG_FEATURE_CHECK_UNICODE_IN_ENV is not set
CONFIG_SUBST_WCHAR=0
CONFIG_LAST_SUPPORTED_WCHAR=0
# CONFIG_UNICODE_COMBINING_WCHARS is not set
# CONFIG_UNICODE_WIDE_WCHARS is not set
# CONFIG_UNICODE_BIDI_SUPPORT is not set
# CONFIG_UNICODE_NEUTRAL_TABLE is not set
# CONFIG_UNICODE_PRESERVE_BROKEN is not set
# CONFIG_LOOP_CONFIGURE is not set
# CONFIG_NO_LOOP_CONFIGURE is not set
CONFIG_TRY_LOOP_CONFIGURE=y

#
# Applets
#

#
# Archival Utilities
#
CONFIG_FEATURE_SEAMLESS_XZ=y
CONFIG_FEATURE_SEAMLESS_LZMA=y
CONFIG_FEATURE_SEAMLESS_BZ2=y
CONFIG_FEATURE_SEAMLESS_GZ=y
CONFIG_FEATURE_SEAMLESS_Z=y
CONFIG_AR=y
CONFIG_FEATURE_AR_LONG_FILENAMES=y
CONFIG_FEATURE_AR_CREATE=y
CONFIG_UNCOMPRESS=y
CONFIG_GUNZIP=y
CONFIG_ZCAT=y
CONFIG_FEATURE_GUNZIP_LONG_OPTIONS=y
CONFIG_BUNZIP2=y
CONFIG_BZCAT=y
CONFIG_UNLZMA=y
CONFIG_LZCAT=y
CONFIG_LZMA=y
CONFIG_UNXZ=y
CONFIG_XZCAT=y
CONFIG_XZ=y
CONFIG_BZIP2=y
CONFIG_BZIP2_SMALL=8
CONFIG_FEATURE_BZIP2_DECOMPRESS=y
CONFIG_CPIO=y
CONFIG_FEATURE_CPIO_O=y
CONFIG_FEATURE_CPIO_P=y
CONFIG_FEATURE_CPIO_IGNORE_DEVNO=y
CONFIG_FEATURE_CPIO_RENUMBER_INODES=y
CONFIG_DPKG=y
CONFIG_DPKG_DEB=y
CONFIG_GZIP=y
CONFIG_FEATURE_GZIP_LONG_OPTIONS=y
CONFIG_GZIP_FAST=0
CONFIG_FEATURE_GZIP_LEVELS=y
CONFIG_FEATURE_GZIP_DECOMPRESS=y
CONFIG_LZOP=y
# CONFIG_UNLZOP is not set
# CONFIG_LZOPCAT is not set
CONFIG_LZOP_COMPR_HIGH=y
CONFIG_RPM=y
CONFIG_RPM2CPIO=y
CONFIG_TAR=y
CONFIG_FEATURE_TAR_LONG_OPTIONS=y
CONFIG_FEATURE_TAR_CREATE=y
CONFIG_FEATURE_TAR_AUTODETECT=y
CONFIG_FEATURE_TAR_FROM=y
CONFIG_FEATURE_TAR_OLDGNU_COMPATIBILITY=y
CONFIG_FEATURE_TAR_OLDSUN_COMPATIBILITY=y
CONFIG_FEATURE_TAR_GNU_EXTENSIONS=y
CONFIG_FEATURE_TAR_TO_COMMAND=y
CONFIG_FEATURE_TAR_UNAME_GNAME=y
CONFIG_FEATURE_TAR_NOPRESERVE_TIME=y
# CONFIG_FEATURE_TAR_SELINUX is not set
CONFIG_UNZIP=y
CONFIG_FEATURE_UNZIP_CDF=y
# CONFIG_FEATURE_UNZIP_BZIP2 is not set
# CONFIG_FEATURE_UNZIP_LZMA is not set
# CONFIG_FEATURE_UNZIP_XZ is not set
CONFIG_FEATURE_LZMA_FAST=y

#
# Coreutils
#
CONFIG_FEATURE_VERBOSE=y

#
# Common options for date and touch
#
# CONFIG_FEATURE_TIMEZONE is not set

#
# Common options for cp and mv
#
CONFIG_FEATURE_PRESERVE_HARDLINKS=y

#
# Common options for df, du, ls
#
CONFIG_FEATURE_HUMAN_READABLE=y
CONFIG_BASENAME=y
CONFIG_CAT=y
CONFIG_FEATURE_CATN=y
CONFIG_FEATURE_CATV=y
CONFIG_CHGRP=y
CONFIG_CHMOD=y
CONFIG_CHOWN=y
CONFIG_FEATURE_CHOWN_LONG_OPTIONS=y
CONFIG_CHROOT=y
CONFIG_CKSUM=y
CONFIG_CRC32=y
CONFIG_COMM=y
CONFIG_CP=y
# CONFIG_FEATURE_CP_LONG_OPTIONS is not set
# CONFIG_FEATURE_CP_REFLINK is not set
CONFIG_CUT=y
CONFIG_FEATURE_CUT_REGEX=y
CONFIG_DATE=y
CONFIG_FEATURE_DATE_ISOFMT=y
# CONFIG_FEATURE_DATE_NANO is not set
CONFIG_FEATURE_DATE_COMPAT=y
CONFIG_DD=y
CONFIG_FEATURE_DD_SIGNAL_HANDLING=y
CONFIG_FEATURE_DD_THIRD_STATUS_LINE=y
CONFIG_FEATURE_DD_IBS_OBS=y
CONFIG_FEATURE_DD_STATUS=y
# CONFIG_DF is not set
# CONFIG_FEATURE_DF_FANCY is not set
# CONFIG_FEATURE_SKIP_ROOTFS is not set
CONFIG_DIRNAME=y
CONFIG_DOS2UNIX=y
CONFIG_UNIX2DOS=y
CONFIG_DU=y
CONFIG_FEATURE_DU_DEFAULT_BLOCKSIZE_1K=y
CONFIG_ECHO=y
CONFIG_FEATURE_FANCY_ECHO=y
# CONFIG_ENV is not set
CONFIG_EXPAND=y
CONFIG_UNEXPAND=y
# CONFIG_EXPR is not set
# CONFIG_EXPR_MATH_SUPPORT_64 is not set
CONFIG_FACTOR=y
CONFIG_FALSE=y
CONFIG_FOLD=y
CONFIG_HEAD=y
CONFIG_FEATURE_FANCY_HEAD=y
# CONFIG_HOSTID is not set
# CONFIG_ID is not set
# CONFIG_GROUPS is not set
CONFIG_INSTALL=y
# CONFIG_FEATURE_INSTALL_LONG_OPTIONS is not set
CONFIG_LINK=y
CONFIG_LN=y
# CONFIG_LOGNAME is not set
CONFIG_LS=y
CONFIG_FEATURE_LS_FILETYPES=y
CONFIG_FEATURE_LS_FOLLOWLINKS=y
CONFIG_FEATURE_LS_RECURSIVE=y
CONFIG_FEATURE_LS_WIDTH=y
CONFIG_FEATURE_LS_SORTFILES=y
CONFIG_FEATURE_LS_TIMESTAMPS=y
CONFIG_FEATURE_LS_USERNAME=y
CONFIG_FEATURE_LS_COLOR=y
CONFIG_FEATURE_LS_COLOR_IS_DEFAULT=y
CONFIG_MD5SUM=y
CONFIG_SHA1SUM=y
CONFIG_SHA256SUM=y
CONFIG_SHA512SUM=y
CONFIG_SHA3SUM=y

#
# Common options for md5sum, sha1sum, sha256sum, sha512sum, sha3sum
#
CONFIG_FEATURE_MD5_SHA1_SUM_CHECK=y
CONFIG_MKDIR=y
CONFIG_MKFIFO=y
CONFIG_MKNOD=y
CONFIG_MKTEMP=y
CONFIG_MV=y
CONFIG_NICE=y
CONFIG_NL=y
CONFIG_NOHUP=y
CONFIG_NPROC=y
CONFIG_OD=y
CONFIG_PASTE=y
CONFIG_PRINTENV=y
CONFIG_PRINTF=y
CONFIG_PWD=y
CONFIG_READLINK=y
CONFIG_FEATURE_READLINK_FOLLOW=y
CONFIG_REALPATH=y
CONFIG_RM=y
CONFIG_RMDIR=y
CONFIG_SEQ=y
CONFIG_SHRED=y
CONFIG_SHUF=y
CONFIG_SLEEP=y
CONFIG_FEATURE_FANCY_SLEEP=y
CONFIG_SORT=y
CONFIG_FEATURE_SORT_BIG=y
# CONFIG_FEATURE_SORT_OPTIMIZE_MEMORY is not set
CONFIG_SPLIT=y
CONFIG_FEATURE_SPLIT_FANCY=y
# CONFIG_STAT is not set
# CONFIG_FEATURE_STAT_FORMAT is not set
# CONFIG_FEATURE_STAT_FILESYSTEM is not set
CONFIG_STTY=y
CONFIG_SUM=y
CONFIG_SYNC=y
CONFIG_FEATURE_SYNC_FANCY=y
# CONFIG_FSYNC is not set
CONFIG_TAC=y
CONFIG_TAIL=y
CONFIG_FEATURE_FANCY_TAIL=y
CONFIG_TEE=y
CONFIG_FEATURE_TEE_USE_BLOCK_IO=y
CONFIG_TEST=y
CONFIG_TEST1=y
CONFIG_TEST2=y
CONFIG_FEATURE_TEST_64=y
CONFIG_TIMEOUT=y
CONFIG_TOUCH=y
CONFIG_FEATURE_TOUCH_SUSV3=y
CONFIG_TR=y
CONFIG_FEATURE_TR_CLASSES=y
CONFIG_FEATURE_TR_EQUIV=y
CONFIG_TRUE=y
CONFIG_TRUNCATE=y
CONFIG_TSORT=y
# CONFIG_TTY is not set
CONFIG_UNAME=y
CONFIG_UNAME_OSNAME="GNU/Linux"
CONFIG_BB_ARCH=y
CONFIG_UNIQ=y
CONFIG_UNLINK=y
# CONFIG_USLEEP is not set
CONFIG_UUDECODE=y
CONFIG_BASE32=y
CONFIG_BASE64=y
CONFIG_UUENCODE=y
CONFIG_WC=y
CONFIG_FEATURE_WC_LARGE=y
# CONFIG_WHO is not set
# CONFIG_W is not set
# CONFIG_USERS is not set
CONFIG_WHOAMI=y
CONFIG_YES=y

#
# Console Utilities
#
CONFIG_CHVT=y
CONFIG_CLEAR=y
CONFIG_DEALLOCVT=y
CONFIG_DUMPKMAP=y
CONFIG_FGCONSOLE=y
# CONFIG_KBD_MODE is not set
# CONFIG_LOADFONT is not set
# CONFIG_SETFONT is not set
# CONFIG_FEATURE_SETFONT_TEXTUAL_MAP is not set
CONFIG_DEFAULT_SETFONT_DIR=""
# CONFIG_FEATURE_LOADFONT_PSF2 is not set
# CONFIG_FEATURE_LOADFONT_RAW is not set
CONFIG_LOADKMAP=y
CONFIG_OPENVT=y
CONFIG_RESET=y
CONFIG_RESIZE=y
CONFIG_FEATURE_RESIZE_PRINT=y
CONFIG_SETCONSOLE=y
# CONFIG_FEATURE_SETCONSOLE_LONG_OPTIONS is not set
CONFIG_SETKEYCODES=y
CONFIG_SETLOGCONS=y
CONFIG_SHOWKEY=y

#
# Debian Utilities
#
CONFIG_PIPE_PROGRESS=y
CONFIG_RUN_PARTS=y
CONFIG_FEATURE_RUN_PARTS_LONG_OPTIONS=y
CONFIG_FEATURE_RUN_PARTS_FANCY=y
CONFIG_START_STOP_DAEMON=y
CONFIG_FEATURE_START_STOP_DAEMON_LONG_OPTIONS=y
CONFIG_FEATURE_START_STOP_DAEMON_FANCY=y
CONFIG_WHICH=y

#
# klibc-utils
#
# CONFIG_MINIPS is not set
# CONFIG_NUKE is not set
CONFIG_RESUME=y
CONFIG_RUN_INIT=y

#
# Editors
#
CONFIG_AWK=y
CONFIG_FEATURE_AWK_LIBM=y
CONFIG_FEATURE_AWK_GNU_EXTENSIONS=y
CONFIG_CMP=y
CONFIG_DIFF=y
CONFIG_FEATURE_DIFF_LONG_OPTIONS=y
CONFIG_FEATURE_DIFF_DIR=y
# CONFIG_ED is not set
CONFIG_PATCH=y
CONFIG_SED=y
CONFIG_VI=y
CONFIG_FEATURE_VI_MAX_LEN=4096
CONFIG_FEATURE_VI_8BIT=y
CONFIG_FEATURE_VI_COLON=y
CONFIG_FEATURE_VI_COLON_EXPAND=y
CONFIG_FEATURE_VI_YANKMARK=y
CONFIG_FEATURE_VI_SEARCH=y
# CONFIG_FEATURE_VI_REGEX_SEARCH is not set
CONFIG_FEATURE_VI_USE_SIGNALS=y
CONFIG_FEATURE_VI_DOT_CMD=y
CONFIG_FEATURE_VI_READONLY=y
CONFIG_FEATURE_VI_SETOPTS=y
CONFIG_FEATURE_VI_SET=y
CONFIG_FEATURE_VI_WIN_RESIZE=y
CONFIG_FEATURE_VI_ASK_TERMINAL=y
CONFIG_FEATURE_VI_UNDO=y
CONFIG_FEATURE_VI_UNDO_QUEUE=y
CONFIG_FEATURE_VI_UNDO_QUEUE_MAX=256
CONFIG_FEATURE_VI_VERBOSE_STATUS=y
CONFIG_FEATURE_ALLOW_EXEC=y

#
# Finding Utilities
#
CONFIG_FIND=y
CONFIG_FEATURE_FIND_PRINT0=y
CONFIG_FEATURE_FIND_MTIME=y
CONFIG_FEATURE_FIND_ATIME=y
CONFIG_FEATURE_FIND_CTIME=y
CONFIG_FEATURE_FIND_MMIN=y
CONFIG_FEATURE_FIND_AMIN=y
CONFIG_FEATURE_FIND_CMIN=y
CONFIG_FEATURE_FIND_PERM=y
CONFIG_FEATURE_FIND_TYPE=y
CONFIG_FEATURE_FIND_EXECUTABLE=y
CONFIG_FEATURE_FIND_XDEV=y
CONFIG_FEATURE_FIND_MAXDEPTH=y
CONFIG_FEATURE_FIND_NEWER=y
CONFIG_FEATURE_FIND_INUM=y
CONFIG_FEATURE_FIND_SAMEFILE=y
CONFIG_FEATURE_FIND_EXEC=y
CONFIG_FEATURE_FIND_EXEC_PLUS=y
CONFIG_FEATURE_FIND_USER=y
CONFIG_FEATURE_FIND_GROUP=y
CONFIG_FEATURE_FIND_NOT=y
CONFIG_FEATURE_FIND_DEPTH=y
CONFIG_FEATURE_FIND_PAREN=y
CONFIG_FEATURE_FIND_SIZE=y
CONFIG_FEATURE_FIND_PRUNE=y
CONFIG_FEATURE_FIND_QUIT=y
CONFIG_FEATURE_FIND_DELETE=y
CONFIG_FEATURE_FIND_EMPTY=y
CONFIG_FEATURE_FIND_PATH=y
CONFIG_FEATURE_FIND_REGEX=y
# CONFIG_FEATURE_FIND_CONTEXT is not set
CONFIG_FEATURE_FIND_LINKS=y
CONFIG_GREP=y
CONFIG_EGREP=y
CONFIG_FGREP=y
# CONFIG_FEATURE_GREP_CONTEXT is not set
CONFIG_XARGS=y
CONFIG_FEATURE_XARGS_SUPPORT_CONFIRMATION=y
CONFIG_FEATURE_XARGS_SUPPORT_QUOTES=y
CONFIG_FEATURE_XARGS_SUPPORT_TERMOPT=y
CONFIG_FEATURE_XARGS_SUPPORT_ZERO_TERM=y
CONFIG_FEATURE_XARGS_SUPPORT_REPL_STR=y
CONFIG_FEATURE_XARGS_SUPPORT_PARALLEL=y
CONFIG_FEATURE_XARGS_SUPPORT_ARGS_FILE=y

#
# Init Utilities
#
# CONFIG_BOOTCHARTD is not set
# CONFIG_FEATURE_BOOTCHARTD_BLOATED_HEADER is not set
# CONFIG_FEATURE_BOOTCHARTD_CONFIG_FILE is not set
CONFIG_HALT=y
CONFIG_POWEROFF=y
CONFIG_REBOOT=y
CONFIG_FEATURE_WAIT_FOR_INIT=y
# CONFIG_FEATURE_CALL_TELINIT is not set
CONFIG_TELINIT_PATH=""
CONFIG_INIT=y
CONFIG_LINUXRC=y
CONFIG_FEATURE_USE_INITTAB=y
# CONFIG_FEATURE_KILL_REMOVED is not set
CONFIG_FEATURE_KILL_DELAY=0
CONFIG_FEATURE_INIT_SCTTY=y
CONFIG_FEATURE_INIT_SYSLOG=y
CONFIG_FEATURE_INIT_QUIET=y
CONFIG_FEATURE_INIT_COREDUMPS=y
CONFIG_INIT_TERMINAL_TYPE="linux"
CONFIG_FEATURE_INIT_MODIFY_CMDLINE=y

#
# Login/Password Management Utilities
#
# CONFIG_FEATURE_SHADOWPASSWDS is not set
# CONFIG_USE_BB_PWD_GRP is not set
# CONFIG_USE_BB_SHADOW is not set
# CONFIG_USE_BB_CRYPT is not set
# CONFIG_USE_BB_CRYPT_SHA is not set
# CONFIG_ADD_SHELL is not set
# CONFIG_REMOVE_SHELL is not set
# CONFIG_ADDGROUP is not set
# CONFIG_FEATURE_ADDUSER_TO_GROUP is not set
# CONFIG_ADDUSER is not set
# CONFIG_FEATURE_CHECK_NAMES is not set
CONFIG_LAST_ID=0
CONFIG_FIRST_SYSTEM_ID=0
CONFIG_LAST_SYSTEM_ID=0
# CONFIG_CHPASSWD is not set
CONFIG_FEATURE_DEFAULT_PASSWD_ALGO=""
# CONFIG_CRYPTPW is not set
CONFIG_MKPASSWD=y
# CONFIG_DELUSER is not set
# CONFIG_DELGROUP is not set
# CONFIG_FEATURE_DEL_USER_FROM_GROUP is not set
# CONFIG_GETTY is not set
# CONFIG_LOGIN is not set
# CONFIG_LOGIN_SESSION_AS_CHILD is not set
# CONFIG_LOGIN_SCRIPTS is not set
# CONFIG_FEATURE_NOLOGIN is not set
# CONFIG_FEATURE_SECURETTY is not set
# CONFIG_PASSWD is not set
# CONFIG_FEATURE_PASSWD_WEAK_CHECK is not set
# CONFIG_SU is not set
# CONFIG_FEATURE_SU_SYSLOG is not set
# CONFIG_FEATURE_SU_CHECKS_SHELLS is not set
# CONFIG_FEATURE_SU_BLANK_PW_NEEDS_SECURE_TTY is not set
# CONFIG_SULOGIN is not set
# CONFIG_VLOCK is not set

#
# Linux Ext2 FS Progs
#
CONFIG_CHATTR=y
# CONFIG_FSCK is not set
CONFIG_LSATTR=y
CONFIG_TUNE2FS=y

#
# Linux Module Utilities
#
CONFIG_MODPROBE_SMALL=y
# CONFIG_DEPMOD is not set
# CONFIG_INSMOD is not set
# CONFIG_LSMOD is not set
# CONFIG_FEATURE_LSMOD_PRETTY_2_6_OUTPUT is not set
CONFIG_MODINFO=y
# CONFIG_MODPROBE is not set
# CONFIG_FEATURE_MODPROBE_BLACKLIST is not set
# CONFIG_RMMOD is not set

#
# Options common to multiple modutils
#
# CONFIG_FEATURE_CMDLINE_MODULE_OPTIONS is not set
# CONFIG_FEATURE_MODPROBE_SMALL_CHECK_ALREADY_LOADED is not set
# CONFIG_FEATURE_2_4_MODULES is not set
# CONFIG_FEATURE_INSMOD_VERSION_CHECKING is not set
# CONFIG_FEATURE_INSMOD_KSYMOOPS_SYMBOLS is not set
# CONFIG_FEATURE_INSMOD_LOADINKMEM is not set
# CONFIG_FEATURE_INSMOD_LOAD_MAP is not set
# CONFIG_FEATURE_INSMOD_LOAD_MAP_FULL is not set
# CONFIG_FEATURE_CHECK_TAINTED_MODULE is not set
# CONFIG_FEATURE_INSMOD_TRY_MMAP is not set
# CONFIG_FEATURE_MODUTILS_ALIAS is not set
# CONFIG_FEATURE_MODUTILS_SYMBOLS is not set
CONFIG_DEFAULT_MODULES_DIR="/lib/modules"
CONFIG_DEFAULT_DEPMOD_FILE="modules.dep"

#
# Linux System Utilities
#
# CONFIG_ACPID is not set
# CONFIG_FEATURE_ACPID_COMPAT is not set
CONFIG_BLKDISCARD=y
CONFIG_BLKID=y
# CONFIG_FEATURE_BLKID_TYPE is not set
CONFIG_BLOCKDEV=y
CONFIG_CAL=y
CONFIG_CHRT=y
CONFIG_DMESG=y
CONFIG_FEATURE_DMESG_PRETTY=y
# CONFIG_EJECT is not set
# CONFIG_FEATURE_EJECT_SCSI is not set
CONFIG_FALLOCATE=y
CONFIG_FATATTR=y
CONFIG_FBSET=y
CONFIG_FEATURE_FBSET_FANCY=y
CONFIG_FEATURE_FBSET_READMODE=y
CONFIG_FDFORMAT=y
CONFIG_FDISK=y
CONFIG_FDISK_SUPPORT_LARGE_DISKS=y
CONFIG_FEATURE_FDISK_WRITABLE=y
# CONFIG_FEATURE_AIX_LABEL is not set
# CONFIG_FEATURE_SGI_LABEL is not set
# CONFIG_FEATURE_SUN_LABEL is not set
# CONFIG_FEATURE_OSF_LABEL is not set
# CONFIG_FEATURE_GPT_LABEL is not set
CONFIG_FEATURE_FDISK_ADVANCED=y
CONFIG_FINDFS=y
CONFIG_FLOCK=y
CONFIG_FDFLUSH=y
CONFIG_FREERAMDISK=y
# CONFIG_FSCK_MINIX is not set
CONFIG_FSFREEZE=y
CONFIG_FSTRIM=y
CONFIG_GETOPT=y
CONFIG_FEATURE_GETOPT_LONG=y
CONFIG_HEXDUMP=y
CONFIG_HD=y
CONFIG_XXD=y
# CONFIG_HWCLOCK is not set
# CONFIG_FEATURE_HWCLOCK_ADJTIME_FHS is not set
# CONFIG_IONICE is not set
# CONFIG_IPCRM is not set
# CONFIG_IPCS is not set
# CONFIG_LAST is not set
# CONFIG_FEATURE_LAST_FANCY is not set
CONFIG_LOSETUP=y
CONFIG_LSPCI=y
CONFIG_LSUSB=y
# CONFIG_MDEV is not set
# CONFIG_FEATURE_MDEV_CONF is not set
# CONFIG_FEATURE_MDEV_RENAME is not set
# CONFIG_FEATURE_MDEV_RENAME_REGEXP is not set
# CONFIG_FEATURE_MDEV_EXEC is not set
# CONFIG_FEATURE_MDEV_LOAD_FIRMWARE is not set
# CONFIG_FEATURE_MDEV_DAEMON is not set
CONFIG_MESG=y
CONFIG_FEATURE_MESG_ENABLE_ONLY_GROUP=y
CONFIG_MKE2FS=y
# CONFIG_MKFS_EXT2 is not set
# CONFIG_MKFS_MINIX is not set
# CONFIG_FEATURE_MINIX2 is not set
# CONFIG_MKFS_REISER is not set
CONFIG_MKDOSFS=y
# CONFIG_MKFS_VFAT is not set
CONFIG_MKSWAP=y
CONFIG_FEATURE_MKSWAP_UUID=y
CONFIG_MORE=y
# CONFIG_MOUNT is not set
# CONFIG_FEATURE_MOUNT_FAKE is not set
# CONFIG_FEATURE_MOUNT_VERBOSE is not set
# CONFIG_FEATURE_MOUNT_HELPERS is not set
# CONFIG_FEATURE_MOUNT_LABEL is not set
# CONFIG_FEATURE_MOUNT_NFS is not set
# CONFIG_FEATURE_MOUNT_CIFS is not set
# CONFIG_FEATURE_MOUNT_FLAGS is not set
# CONFIG_FEATURE_MOUNT_FSTAB is not set
# CONFIG_FEATURE_MOUNT_OTHERTAB is not set
# CONFIG_MOUNTPOINT is not set
CONFIG_NOLOGIN=y
# CONFIG_NOLOGIN_DEPENDENCIES is not set
CONFIG_NSENTER=y
# CONFIG_PIVOT_ROOT is not set
# CONFIG_RDATE is not set
CONFIG_RDEV=y
CONFIG_READPROFILE=y
CONFIG_RENICE=y
CONFIG_REV=y
CONFIG_RTCWAKE=y
CONFIG_SCRIPT=y
CONFIG_SCRIPTREPLAY=y
# CONFIG_SETARCH is not set
CONFIG_LINUX32=y
CONFIG_LINUX64=y
CONFIG_SETPRIV=y
CONFIG_FEATURE_SETPRIV_DUMP=y
CONFIG_FEATURE_SETPRIV_CAPABILITIES=y
CONFIG_FEATURE_SETPRIV_CAPABILITY_NAMES=y
CONFIG_SETSID=y
# CONFIG_SWAPON is not set
# CONFIG_FEATURE_SWAPON_DISCARD is not set
# CONFIG_FEATURE_SWAPON_PRI is not set
# CONFIG_SWAPOFF is not set
# CONFIG_FEATURE_SWAPONOFF_LABEL is not set
# CONFIG_SWITCH_ROOT is not set
# CONFIG_TASKSET is not set
# CONFIG_FEATURE_TASKSET_FANCY is not set
# CONFIG_FEATURE_TASKSET_CPULIST is not set
CONFIG_UEVENT=y
# CONFIG_UMOUNT is not set
# CONFIG_FEATURE_UMOUNT_ALL is not set
CONFIG_UNSHARE=y
# CONFIG_WALL is not set
# CONFIG_FEATURE_MOUNT_LOOP is not set
# CONFIG_FEATURE_MOUNT_LOOP_CREATE is not set
# CONFIG_FEATURE_MTAB_SUPPORT is not set
CONFIG_VOLUMEID=y

#
# Filesystem/Volume identification
#
CONFIG_FEATURE_VOLUMEID_BCACHE=y
CONFIG_FEATURE_VOLUMEID_BTRFS=y
CONFIG_FEATURE_VOLUMEID_CRAMFS=y
CONFIG_FEATURE_VOLUMEID_EROFS=y
CONFIG_FEATURE_VOLUMEID_EXFAT=y
CONFIG_FEATURE_VOLUMEID_EXT=y
CONFIG_FEATURE_VOLUMEID_F2FS=y
CONFIG_FEATURE_VOLUMEID_FAT=y
CONFIG_FEATURE_VOLUMEID_HFS=y
CONFIG_FEATURE_VOLUMEID_ISO9660=y
CONFIG_FEATURE_VOLUMEID_JFS=y
# CONFIG_FEATURE_VOLUMEID_LFS is not set
CONFIG_FEATURE_VOLUMEID_LINUXRAID=y
CONFIG_FEATURE_VOLUMEID_LINUXSWAP=y
CONFIG_FEATURE_VOLUMEID_LUKS=y
CONFIG_FEATURE_VOLUMEID_MINIX=y
CONFIG_FEATURE_VOLUMEID_NILFS=y
CONFIG_FEATURE_VOLUMEID_NTFS=y
CONFIG_FEATURE_VOLUMEID_OCFS2=y
CONFIG_FEATURE_VOLUMEID_REISERFS=y
CONFIG_FEATURE_VOLUMEID_ROMFS=y
# CONFIG_FEATURE_VOLUMEID_SQUASHFS is not set
CONFIG_FEATURE_VOLUMEID_SYSV=y
CONFIG_FEATURE_VOLUMEID_UBIFS=y
CONFIG_FEATURE_VOLUMEID_UDF=y
CONFIG_FEATURE_VOLUMEID_XFS=y

#
# Miscellaneous Utilities
#
# CONFIG_ADJTIMEX is not set
CONFIG_ASCII=y
# CONFIG_BBCONFIG is not set
# CONFIG_FEATURE_COMPRESS_BBCONFIG is not set
CONFIG_BC=y
CONFIG_DC=y
CONFIG_FEATURE_DC_BIG=y
# CONFIG_FEATURE_DC_LIBM is not set
CONFIG_FEATURE_BC_INTERACTIVE=y
CONFIG_FEATURE_BC_LONG_OPTIONS=y
CONFIG_BEEP=y
CONFIG_FEATURE_BEEP_FREQ=4000
CONFIG_FEATURE_BEEP_LENGTH_MS=30
CONFIG_CHAT=y
CONFIG_FEATURE_CHAT_NOFAIL=y
# CONFIG_FEATURE_CHAT_TTY_HIFI is not set
CONFIG_FEATURE_CHAT_IMPLICIT_CR=y
CONFIG_FEATURE_CHAT_SWALLOW_OPTS=y
CONFIG_FEATURE_CHAT_SEND_ESCAPES=y
CONFIG_FEATURE_CHAT_VAR_ABORT_LEN=y
CONFIG_FEATURE_CHAT_CLR_ABORT=y
# CONFIG_CONSPY is not set
# CONFIG_CROND is not set
# CONFIG_FEATURE_CROND_D is not set
# CONFIG_FEATURE_CROND_CALL_SENDMAIL is not set
# CONFIG_FEATURE_CROND_SPECIAL_TIMES is not set
CONFIG_FEATURE_CROND_DIR=""
# CONFIG_CRONTAB is not set
# CONFIG_DEVFSD is not set
# CONFIG_DEVFSD_MODLOAD is not set
# CONFIG_DEVFSD_FG_NP is not set
# CONFIG_DEVFSD_VERBOSE is not set
# CONFIG_FEATURE_DEVFS is not set
CONFIG_DEVMEM=y
CONFIG_FBSPLASH=y
# CONFIG_FLASH_ERASEALL is not set
CONFIG_FLASH_LOCK=y
CONFIG_FLASH_UNLOCK=y
CONFIG_FLASHCP=y
CONFIG_HDPARM=y
CONFIG_FEATURE_HDPARM_GET_IDENTITY=y
CONFIG_FEATURE_HDPARM_HDIO_SCAN_HWIF=y
CONFIG_FEATURE_HDPARM_HDIO_UNREGISTER_HWIF=y
CONFIG_FEATURE_HDPARM_HDIO_DRIVE_RESET=y
CONFIG_FEATURE_HDPARM_HDIO_TRISTATE_HWIF=y
CONFIG_FEATURE_HDPARM_HDIO_GETSET_DMA=y
CONFIG_HEXEDIT=y
CONFIG_I2CGET=y
CONFIG_I2CSET=y
CONFIG_I2CDUMP=y
CONFIG_I2CDETECT=y
CONFIG_I2CTRANSFER=y
CONFIG_INOTIFYD=y
# CONFIG_LESS is not set
CONFIG_FEATURE_LESS_MAXLINES=0
# CONFIG_FEATURE_LESS_BRACKETS is not set
# CONFIG_FEATURE_LESS_FLAGS is not set
# CONFIG_FEATURE_LESS_TRUNCATE is not set
# CONFIG_FEATURE_LESS_MARKS is not set
# CONFIG_FEATURE_LESS_REGEXP is not set
# CONFIG_FEATURE_LESS_WINCH is not set
# CONFIG_FEATURE_LESS_ASK_TERMINAL is not set
# CONFIG_FEATURE_LESS_DASHCMD is not set
# CONFIG_FEATURE_LESS_LINENUMS is not set
# CONFIG_FEATURE_LESS_RAW is not set
# CONFIG_FEATURE_LESS_ENV is not set
CONFIG_LSSCSI=y
CONFIG_MAKEDEVS=y
# CONFIG_FEATURE_MAKEDEVS_LEAF is not set
CONFIG_FEATURE_MAKEDEVS_TABLE=y
CONFIG_MAN=y
# CONFIG_MICROCOM is not set
CONFIG_MIM=y
# CONFIG_MT is not set
# CONFIG_NANDWRITE is not set
CONFIG_NANDDUMP=y
CONFIG_PARTPROBE=y
CONFIG_RAIDAUTORUN=y
# CONFIG_READAHEAD is not set
# CONFIG_RFKILL is not set
# CONFIG_RUNLEVEL is not set
CONFIG_RX=y
CONFIG_SEEDRNG=y
CONFIG_SETFATTR=y
CONFIG_SETSERIAL=y
CONFIG_STRINGS=y
CONFIG_TIME=y
CONFIG_TREE=y
CONFIG_TS=y
CONFIG_TTYSIZE=y
# CONFIG_UBIATTACH is not set
# CONFIG_UBIDETACH is not set
# CONFIG_UBIMKVOL is not set
# CONFIG_UBIRMVOL is not set
# CONFIG_UBIRSVOL is not set
# CONFIG_UBIUPDATEVOL is not set
CONFIG_UBIRENAME=y
CONFIG_VOLNAME=y
# CONFIG_WATCHDOG is not set
# CONFIG_FEATURE_WATCHDOG_OPEN_TWICE is not set

#
# Networking Utilities
#
# CONFIG_FEATURE_IPV6 is not set
# CONFIG_FEATURE_UNIX_LOCAL is not set
# CONFIG_FEATURE_PREFER_IPV4_ADDRESS is not set
CONFIG_VERBOSE_RESOLUTION_ERRORS=y
# CONFIG_FEATURE_ETC_NETWORKS is not set
# CONFIG_FEATURE_ETC_SERVICES is not set
# CONFIG_FEATURE_HWIB is not set
# CONFIG_FEATURE_TLS_SHA1 is not set
CONFIG_ARP=y
# CONFIG_ARPING is not set
# CONFIG_BRCTL is not set
# CONFIG_FEATURE_BRCTL_FANCY is not set
# CONFIG_FEATURE_BRCTL_SHOW is not set
CONFIG_DNSD=y
# CONFIG_ETHER_WAKE is not set
CONFIG_FTPD=y
CONFIG_FEATURE_FTPD_WRITE=y
CONFIG_FEATURE_FTPD_ACCEPT_BROKEN_LIST=y
CONFIG_FEATURE_FTPD_AUTHENTICATION=y
CONFIG_FTPGET=y
CONFIG_FTPPUT=y
# CONFIG_FEATURE_FTPGETPUT_LONG_OPTIONS is not set
# CONFIG_HOSTNAME is not set
CONFIG_DNSDOMAINNAME=y
CONFIG_HTTPD=y
CONFIG_FEATURE_HTTPD_PORT_DEFAULT=80
CONFIG_FEATURE_HTTPD_RANGES=y
CONFIG_FEATURE_HTTPD_SETUID=y
CONFIG_FEATURE_HTTPD_BASIC_AUTH=y
# CONFIG_FEATURE_HTTPD_AUTH_MD5 is not set
CONFIG_FEATURE_HTTPD_CGI=y
CONFIG_FEATURE_HTTPD_CONFIG_WITH_SCRIPT_INTERPR=y
CONFIG_FEATURE_HTTPD_SET_REMOTE_PORT_TO_ENV=y
CONFIG_FEATURE_HTTPD_ENCODE_URL_STR=y
CONFIG_FEATURE_HTTPD_ERROR_PAGES=y
CONFIG_FEATURE_HTTPD_PROXY=y
CONFIG_FEATURE_HTTPD_GZIP=y
CONFIG_FEATURE_HTTPD_ETAG=y
CONFIG_FEATURE_HTTPD_LAST_MODIFIED=y
CONFIG_FEATURE_HTTPD_DATE=y
CONFIG_FEATURE_HTTPD_ACL_IP=y
CONFIG_IFCONFIG=y
CONFIG_FEATURE_IFCONFIG_STATUS=y
# CONFIG_FEATURE_IFCONFIG_SLIP is not set
CONFIG_FEATURE_IFCONFIG_MEMSTART_IOADDR_IRQ=y
CONFIG_FEATURE_IFCONFIG_HW=y
CONFIG_FEATURE_IFCONFIG_BROADCAST_PLUS=y
# CONFIG_IFENSLAVE is not set
# CONFIG_IFPLUGD is not set
CONFIG_IFUP=y
CONFIG_IFDOWN=y
CONFIG_IFUPDOWN_IFSTATE_PATH="/var/run/ifstate"
CONFIG_FEATURE_IFUPDOWN_IP=y
CONFIG_FEATURE_IFUPDOWN_IPV4=y
# CONFIG_FEATURE_IFUPDOWN_IPV6 is not set
CONFIG_FEATURE_IFUPDOWN_MAPPING=y
# CONFIG_FEATURE_IFUPDOWN_EXTERNAL_DHCP is not set
# CONFIG_INETD is not set
# CONFIG_FEATURE_INETD_SUPPORT_BUILTIN_ECHO is not set
# CONFIG_FEATURE_INETD_SUPPORT_BUILTIN_DISCARD is not set
# CONFIG_FEATURE_INETD_SUPPORT_BUILTIN_TIME is not set
# CONFIG_FEATURE_INETD_SUPPORT_BUILTIN_DAYTIME is not set
# CONFIG_FEATURE_INETD_SUPPORT_BUILTIN_CHARGEN is not set
# CONFIG_FEATURE_INETD_RPC is not set
CONFIG_IP=y
CONFIG_IPADDR=y
CONFIG_IPLINK=y
CONFIG_IPROUTE=y
CONFIG_IPTUNNEL=y
CONFIG_IPRULE=y
CONFIG_IPNEIGH=y
CONFIG_FEATURE_IP_ADDRESS=y
CONFIG_FEATURE_IP_LINK=y
CONFIG_FEATURE_IP_ROUTE=y
CONFIG_FEATURE_IP_ROUTE_DIR="/etc/iproute2"
CONFIG_FEATURE_IP_TUNNEL=y
CONFIG_FEATURE_IP_RULE=y
CONFIG_FEATURE_IP_NEIGH=y
# CONFIG_FEATURE_IP_RARE_PROTOCOLS is not set
CONFIG_IPCALC=y
# CONFIG_FEATURE_IPCALC_LONG_OPTIONS is not set
CONFIG_FEATURE_IPCALC_FANCY=y
CONFIG_FAKEIDENTD=y
# CONFIG_NAMEIF is not set
# CONFIG_FEATURE_NAMEIF_EXTENDED is not set
CONFIG_NBDCLIENT=y
CONFIG_NC=y
# CONFIG_NETCAT is not set
CONFIG_NC_SERVER=y
CONFIG_NC_EXTRA=y
# CONFIG_NC_110_COMPAT is not set
CONFIG_NETSTAT=y
CONFIG_FEATURE_NETSTAT_WIDE=y
CONFIG_FEATURE_NETSTAT_PRG=y
CONFIG_NSLOOKUP=y
# CONFIG_FEATURE_NSLOOKUP_BIG is not set
# CONFIG_FEATURE_NSLOOKUP_LONG_OPTIONS is not set
# CONFIG_NTPD is not set
# CONFIG_FEATURE_NTPD_SERVER is not set
# CONFIG_FEATURE_NTPD_CONF is not set
# CONFIG_FEATURE_NTP_AUTH is not set
# CONFIG_PING is not set
# CONFIG_PING6 is not set
# CONFIG_FEATURE_FANCY_PING is not set
CONFIG_PSCAN=y
CONFIG_ROUTE=y
# CONFIG_SLATTACH is not set
CONFIG_SSL_CLIENT=y
CONFIG_TC=y
CONFIG_FEATURE_TC_INGRESS=y
CONFIG_TCPSVD=y
# CONFIG_UDPSVD is not set
# CONFIG_TELNET is not set
# CONFIG_FEATURE_TELNET_TTYPE is not set
# CONFIG_FEATURE_TELNET_AUTOLOGIN is not set
# CONFIG_FEATURE_TELNET_WIDTH is not set
# CONFIG_TELNETD is not set
# CONFIG_FEATURE_TELNETD_STANDALONE is not set
CONFIG_FEATURE_TELNETD_PORT_DEFAULT=0
# CONFIG_FEATURE_TELNETD_INETD_WAIT is not set
# CONFIG_TFTP is not set
# CONFIG_FEATURE_TFTP_PROGRESS_BAR is not set
# CONFIG_FEATURE_TFTP_HPA_COMPAT is not set
# CONFIG_TFTPD is not set
# CONFIG_FEATURE_TFTP_GET is not set
# CONFIG_FEATURE_TFTP_PUT is not set
# CONFIG_FEATURE_TFTP_BLOCKSIZE is not set
# CONFIG_TFTP_DEBUG is not set
CONFIG_TLS=y
# CONFIG_TRACEROUTE is not set
# CONFIG_TRACEROUTE6 is not set
# CONFIG_FEATURE_TRACEROUTE_VERBOSE is not set
# CONFIG_FEATURE_TRACEROUTE_USE_ICMP is not set
CONFIG_TUNCTL=y
CONFIG_FEATURE_TUNCTL_UG=y
# CONFIG_VCONFIG is not set
CONFIG_WGET=y
CONFIG_FEATURE_WGET_LONG_OPTIONS=y
CONFIG_FEATURE_WGET_STATUSBAR=y
CONFIG_FEATURE_WGET_FTP=y
CONFIG_FEATURE_WGET_AUTHENTICATION=y
CONFIG_FEATURE_WGET_TIMEOUT=y
CONFIG_FEATURE_WGET_HTTPS=y
CONFIG_FEATURE_WGET_OPENSSL=y
CONFIG_WHOIS=y
# CONFIG_ZCIP is not set
# CONFIG_UDHCPD is not set
# CONFIG_FEATURE_UDHCPD_BASE_IP_ON_MAC is not set
# CONFIG_FEATURE_UDHCPD_WRITE_LEASES_EARLY is not set
CONFIG_DHCPD_LEASES_FILE=""
# CONFIG_DUMPLEASES is not set
# CONFIG_DHCPRELAY is not set
CONFIG_UDHCPC=y
CONFIG_FEATURE_UDHCPC_ARPING=y
CONFIG_FEATURE_UDHCPC_SANITIZEOPT=y
CONFIG_UDHCPC_DEFAULT_SCRIPT="/usr/share/udhcpc/default.script"
CONFIG_UDHCPC6_DEFAULT_SCRIPT=""
# CONFIG_UDHCPC6 is not set
# CONFIG_FEATURE_UDHCPC6_RFC3646 is not set
# CONFIG_FEATURE_UDHCPC6_RFC4704 is not set
# CONFIG_FEATURE_UDHCPC6_RFC4833 is not set
# CONFIG_FEATURE_UDHCPC6_RFC5970 is not set

#
# Common options for DHCP applets
#
CONFIG_UDHCPC_DEFAULT_INTERFACE="eth0"
# CONFIG_FEATURE_UDHCP_PORT is not set
CONFIG_UDHCP_DEBUG=9
CONFIG_UDHCPC_SLACK_FOR_BUGGY_SERVERS=80
CONFIG_FEATURE_UDHCP_RFC3397=y
CONFIG_FEATURE_UDHCP_8021Q=y
CONFIG_IFUPDOWN_UDHCPC_CMD_OPTIONS="-R -n"

#
# Print Utilities
#
CONFIG_LPD=y
CONFIG_LPR=y
CONFIG_LPQ=y

#
# Mail Utilities
#
CONFIG_FEATURE_MIME_CHARSET="us-ascii"
CONFIG_MAKEMIME=y
CONFIG_POPMAILDIR=y
CONFIG_FEATURE_POPMAILDIR_DELIVERY=y
CONFIG_REFORMIME=y
CONFIG_FEATURE_REFORMIME_COMPAT=y
CONFIG_SENDMAIL=y

#
# Process Utilities
#
# CONFIG_FEATURE_FAST_TOP is not set
CONFIG_FEATURE_SHOW_THREADS=y
# CONFIG_FREE is not set
CONFIG_FUSER=y
CONFIG_IOSTAT=y
# CONFIG_KILL is not set
# CONFIG_KILLALL is not set
# CONFIG_KILLALL5 is not set
CONFIG_LSOF=y
CONFIG_MPSTAT=y
CONFIG_NMETER=y
# CONFIG_PGREP is not set
# CONFIG_PKILL is not set
CONFIG_PIDOF=y
CONFIG_FEATURE_PIDOF_SINGLE=y
CONFIG_FEATURE_PIDOF_OMIT=y
CONFIG_PMAP=y
CONFIG_POWERTOP=y
CONFIG_FEATURE_POWERTOP_INTERACTIVE=y
# CONFIG_PS is not set
# CONFIG_FEATURE_PS_WIDE is not set
# CONFIG_FEATURE_PS_LONG is not set
# CONFIG_FEATURE_PS_TIME is not set
# CONFIG_FEATURE_PS_UNUSUAL_SYSTEMS is not set
# CONFIG_FEATURE_PS_ADDITIONAL_COLUMNS is not set
CONFIG_PSTREE=y
CONFIG_PWDX=y
CONFIG_SMEMCAP=y
CONFIG_BB_SYSCTL=y
CONFIG_TOP=y
CONFIG_FEATURE_TOP_INTERACTIVE=y
CONFIG_FEATURE_TOP_CPU_USAGE_PERCENTAGE=y
CONFIG_FEATURE_TOP_CPU_GLOBAL_PERCENTS=y
CONFIG_FEATURE_TOP_SMP_CPU=y
CONFIG_FEATURE_TOP_DECIMALS=y
CONFIG_FEATURE_TOP_SMP_PROCESS=y
CONFIG_FEATURE_TOPMEM=y
# CONFIG_UPTIME is not set
# CONFIG_FEATURE_UPTIME_UTMP_SUPPORT is not set
CONFIG_WATCH=y

#
# Runit Utilities
#
CONFIG_CHPST=y
CONFIG_SETUIDGID=y
CONFIG_ENVUIDGID=y
CONFIG_ENVDIR=y
CONFIG_SOFTLIMIT=y
CONFIG_RUNSV=y
CONFIG_RUNSVDIR=y
# CONFIG_FEATURE_RUNSVDIR_LOG is not set
CONFIG_SV=y
CONFIG_SV_DEFAULT_SERVICE_DIR="/var/service"
CONFIG_SVC=y
CONFIG_SVOK=y
CONFIG_SVLOGD=y
# CONFIG_CHCON is not set
# CONFIG_GETENFORCE is not set
# CONFIG_GETSEBOOL is not set
# CONFIG_LOAD_POLICY is not set
# CONFIG_MATCHPATHCON is not set
# CONFIG_RUNCON is not set
# CONFIG_SELINUXENABLED is not set
# CONFIG_SESTATUS is not set
# CONFIG_SETENFORCE is not set
# CONFIG_SETFILES is not set
# CONFIG_FEATURE_SETFILES_CHECK_OPTION is not set
# CONFIG_RESTORECON is not set
# CONFIG_SETSEBOOL is not set

#
# Shells
#
CONFIG_SH_IS_ASH=y
# CONFIG_SH_IS_HUSH is not set
# CONFIG_SH_IS_NONE is not set
# CONFIG_BASH_IS_ASH is not set
# CONFIG_BASH_IS_HUSH is not set
CONFIG_BASH_IS_NONE=y
CONFIG_SHELL_ASH=y
CONFIG_ASH=y
# CONFIG_ASH_OPTIMIZE_FOR_SIZE is not set
CONFIG_ASH_INTERNAL_GLOB=y
CONFIG_ASH_BASH_COMPAT=y
CONFIG_ASH_BASH_SOURCE_CURDIR=y
CONFIG_ASH_BASH_NOT_FOUND_HOOK=y
CONFIG_ASH_JOB_CONTROL=y
CONFIG_ASH_ALIAS=y
CONFIG_ASH_RANDOM_SUPPORT=y
CONFIG_ASH_EXPAND_PRMT=y
# CONFIG_ASH_IDLE_TIMEOUT is not set
# CONFIG_ASH_MAIL is not set
CONFIG_ASH_ECHO=y
CONFIG_ASH_PRINTF=y
CONFIG_ASH_TEST=y
CONFIG_ASH_SLEEP=y
CONFIG_ASH_HELP=y
CONFIG_ASH_GETOPTS=y
CONFIG_ASH_CMDCMD=y
CONFIG_CTTYHACK=y
# CONFIG_HUSH is not set
CONFIG_SHELL_HUSH=y
CONFIG_HUSH_BASH_COMPAT=y
CONFIG_HUSH_BRACE_EXPANSION=y
# CONFIG_HUSH_BASH_SOURCE_CURDIR is not set
CONFIG_HUSH_LINENO_VAR=y
CONFIG_HUSH_INTERACTIVE=y
CONFIG_HUSH_SAVEHISTORY=y
CONFIG_HUSH_JOB=y
CONFIG_HUSH_TICK=y
CONFIG_HUSH_IF=y
CONFIG_HUSH_LOOPS=y
CONFIG_HUSH_CASE=y
CONFIG_HUSH_FUNCTIONS=y
CONFIG_HUSH_LOCAL=y
CONFIG_HUSH_RANDOM_SUPPORT=y
CONFIG_HUSH_MODE_X=y
CONFIG_HUSH_ECHO=y
CONFIG_HUSH_PRINTF=y
CONFIG_HUSH_TEST=y
CONFIG_HUSH_HELP=y
CONFIG_HUSH_EXPORT=y
CONFIG_HUSH_EXPORT_N=y
CONFIG_HUSH_READONLY=y
CONFIG_HUSH_KILL=y
CONFIG_HUSH_WAIT=y
CONFIG_HUSH_COMMAND=y
CONFIG_HUSH_TRAP=y
CONFIG_HUSH_TYPE=y
CONFIG_HUSH_TIMES=y
CONFIG_HUSH_READ=y
CONFIG_HUSH_SET=y
CONFIG_HUSH_UNSET=y
CONFIG_HUSH_ULIMIT=y
CONFIG_HUSH_UMASK=y
CONFIG_HUSH_GETOPTS=y
# CONFIG_HUSH_MEMLEAK is not set

#
# Options common to all shells
#
CONFIG_FEATURE_SH_MATH=y
CONFIG_FEATURE_SH_MATH_64=y
CONFIG_FEATURE_SH_MATH_BASE=y
# CONFIG_FEATURE_SH_EXTRA_QUIET is not set
CONFIG_FEATURE_SH_STANDALONE=y
CONFIG_FEATURE_SH_NOFORK=y
CONFIG_FEATURE_SH_READ_FRAC=y
# CONFIG_FEATURE_SH_HISTFILESIZE is not set
CONFIG_FEATURE_SH_EMBEDDED_SCRIPTS=y

#
# System Logging Utilities
#
CONFIG_KLOGD=y
CONFIG_FEATURE_KLOGD_KLOGCTL=y
# CONFIG_LOGGER is not set
# CONFIG_LOGREAD is not set
# CONFIG_FEATURE_LOGREAD_REDUCED_LOCKING is not set
# CONFIG_SYSLOGD is not set
# CONFIG_FEATURE_ROTATE_LOGFILE is not set
# CONFIG_FEATURE_REMOTE_LOG is not set
# CONFIG_FEATURE_SYSLOGD_DUP is not set
# CONFIG_FEATURE_SYSLOGD_CFG is not set
# CONFIG_FEATURE_SYSLOGD_PRECISE_TIMESTAMPS is not set
CONFIG_FEATURE_SYSLOGD_READ_BUFFER_SIZE=0
# CONFIG_FEATURE_IPC_SYSLOG is not set
CONFIG_FEATURE_IPC_SYSLOG_BUFFER_SIZE=0
# CONFIG_FEATURE_KMSG_SYSLOG is not set

#
# dowork
#
CONFIG_DOWORK=y
